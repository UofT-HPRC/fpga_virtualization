`timescale 1ns / 1ps
`default_nettype none

/*
Shell Wrapper for physical layer interfaces (for the Alveo U200 platform)

Author: Daniel Rozhko, PhD Candidate University of Toronto

Description:
   This module wraps all of the physcial layer interfaces needed by the
   shell, which includes a network interface (TX and RX) and some control 
   interface (e.g. PCIe).

Parameters:
   NET_AXIS_BUS_WIDTH - the data width of the axi-streams (must be multiple of 8)
   NET_MAX_PACKET_LENGTH - the maximum network packet length to support (for forced tlast)

Ports:
   axis_tx_s_* - the input axi stream for the tx direction, to phy
   axis_rx_m_* - the output axi stream for the rx direction, from phy
   axis_aclk - clock to which all of the network signals are synchronous (generated by physical layer)
   axis_aresetn - active-low reset corresponding to above clock (generated by physical layer)

   top_ctrl_* - the AXI-Lite control interface for the top-level control (e.g. PCIe)
   top_mem_* - the AXI4 memory-access interface for the top-level (e.g. PCIe)
   top_aclk - clock to which the control signal is synchronous (generated by physical layer)
   top_aresetn - active-low reset corresponding to above clock (generated by physical layer)

*/


module phy_shell
#(
    //Network AXI Stream Params (as seen by application regions)
    parameter NET_AXIS_BUS_WIDTH = 64,

    //Network Packet Params
    parameter NET_MAX_PACKET_LENGTH = 1522



    //AXI-Lite Interface Params
    //parameter CTRL_AXI_DATA_WIDTH = 32, //Fixed to 32 for now, 64-bit not supported by some cores
)
(
    //Egress Output AXI stream (TX packets to Phy)
    input wire [NET_AXIS_BUS_WIDTH-1:0]          axis_tx_0_s_tdata,
    input wire [(NET_AXIS_BUS_WIDTH/8)-1:0]      axis_tx_0_s_tkeep,
    input wire                                   axis_tx_0_s_tlast,
    input wire                                   axis_tx_0_s_tvalid,
    output wire                                  axis_tx_0_s_tready,

    //Ingress Input AXI stream (RX packets from Phy)
    output wire [NET_AXIS_BUS_WIDTH-1:0]         axis_rx_0_m_tdata,
    output wire [(NET_AXIS_BUS_WIDTH/8)-1:0]     axis_rx_0_m_tkeep,
    output wire                                  axis_rx_0_m_tlast,
    output wire                                  axis_rx_0_m_tvalid,
    input wire                                   axis_rx_0_m_tready,

    //Egress Output AXI stream (TX packets to Phy)
    input wire [NET_AXIS_BUS_WIDTH-1:0]          axis_tx_1_s_tdata,
    input wire [(NET_AXIS_BUS_WIDTH/8)-1:0]      axis_tx_1_s_tkeep,
    input wire                                   axis_tx_1_s_tlast,
    input wire                                   axis_tx_1_s_tvalid,
    output wire                                  axis_tx_1_s_tready,

    //Ingress Input AXI stream (RX packets from Phy)
    output wire [NET_AXIS_BUS_WIDTH-1:0]         axis_rx_1_m_tdata,
    output wire [(NET_AXIS_BUS_WIDTH/8)-1:0]     axis_rx_1_m_tkeep,
    output wire                                  axis_rx_1_m_tlast,
    output wire                                  axis_rx_1_m_tvalid,
    input wire                                   axis_rx_1_m_tready,

    //Network Clocking
    output wire  axis_aclk,
    output wire  axis_aresetn,
    


    //The AXI-Lite Control Interface (from control, e.g. PCIe)
    //Write Address Channel  
    output wire  [31:0]                        top_ctrl_awaddr,
    output wire                                top_ctrl_awvalid,
    input wire                                 top_ctrl_awready,
    //Write Data Channel
    output wire  [31:0]                        top_ctrl_wdata,
    output wire  [3:0]                         top_ctrl_wstrb,
    output wire                                top_ctrl_wvalid,
    input wire                                 top_ctrl_wready,
    //Write Response Channel
    input wire [1:0]                           top_ctrl_bresp,
    input wire                                 top_ctrl_bvalid,
    output wire                                top_ctrl_bready,
    //Read Address Channel 
    output wire  [31:0]                        top_ctrl_araddr,
    output wire                                top_ctrl_arvalid,
    input wire                                 top_ctrl_arready,
    //Read Data Response Channel
    input wire [31:0]                          top_ctrl_rdata,
    input wire [1:0]                           top_ctrl_rresp,
    input wire                                 top_ctrl_rvalid,
    output wire                                top_ctrl_rready,

    //Ctrl Clocking
    output wire  top_aclk,
    output wire  top_aresetn,
    
    //Physical layer ports (from include file)
    `include "phy_signals.svh"
);

    //--------------------------------------------------------//
    //   PHY layer defined in BD                              //
    //--------------------------------------------------------//

    //TODO - update this
    phy_bd_wrapper phy_bd_inst
    (
        .M_AXI_LITE_araddr  (top_ctrl_araddr),
        .M_AXI_LITE_arprot  ( ),
        .M_AXI_LITE_arready (top_ctrl_arready),
        .M_AXI_LITE_arvalid (top_ctrl_arvalid),
        .M_AXI_LITE_awaddr  (top_ctrl_awaddr),
        .M_AXI_LITE_awprot  ( ),
        .M_AXI_LITE_awready (top_ctrl_awready),
        .M_AXI_LITE_awvalid (top_ctrl_awvalid),
        .M_AXI_LITE_bready  (top_ctrl_bready),
        .M_AXI_LITE_bresp   (top_ctrl_bresp),
        .M_AXI_LITE_bvalid  (top_ctrl_bvalid),
        .M_AXI_LITE_rdata   (top_ctrl_rdata),
        .M_AXI_LITE_rready  (top_ctrl_rready),
        .M_AXI_LITE_rresp   (top_ctrl_rresp),
        .M_AXI_LITE_rvalid  (top_ctrl_rvalid),
        .M_AXI_LITE_wdata   (top_ctrl_wdata),
        .M_AXI_LITE_wready  (top_ctrl_wready),
        .M_AXI_LITE_wstrb   (top_ctrl_wstrb),
        .M_AXI_LITE_wvalid  (top_ctrl_wvalid),
        
        .pcie_aclk          (top_aclk),
        .pcie_aresetn       (top_aresetn),
    
        .axis_rx_tdata      (axis_rx_0_m_tdata),
        .axis_rx_tkeep      (axis_rx_0_m_tkeep),
        .axis_rx_tlast      (axis_rx_0_m_tlast),
        .axis_rx_tuser      ( ),
        .axis_rx_tvalid     (axis_rx_0_m_tvalid),
    
        .axis_tx_tdata      (axis_tx_0_s_tdata),
        .axis_tx_tkeep      (axis_tx_0_s_tkeep),
        .axis_tx_tlast      (axis_tx_0_s_tlast),
        .axis_tx_tready     (axis_tx_0_s_tready),
        .axis_tx_tuser      (1'b0),
        .axis_tx_tvalid     (axis_tx_0_s_tvalid),

        .axis_rx_tdata      (axis_rx_1_m_tdata),
        .axis_rx_tkeep      (axis_rx_1_m_tkeep),
        .axis_rx_tlast      (axis_rx_1_m_tlast),
        .axis_rx_tuser      ( ),
        .axis_rx_tvalid     (axis_rx_1_m_tvalid),
    
        .axis_tx_tdata      (axis_tx_1_s_tdata),
        .axis_tx_tkeep      (axis_tx_1_s_tkeep),
        .axis_tx_tlast      (axis_tx_1_s_tlast),
        .axis_tx_tready     (axis_tx_1_s_tready),
        .axis_tx_tuser      (1'b0),
        .axis_tx_tvalid     (axis_tx_1_s_tvalid),
        
        .qsfp0_aclk         (axis_aclk),
        .qsfp0_aresetn      (axis_aresetn),
    
        .pci_express_x1_rxn  (pci_express_x1_rxn),
        .pci_express_x1_rxp  (pci_express_x1_rxp),
        .pci_express_x1_txn  (pci_express_x1_txn),
        .pci_express_x1_txp  (pci_express_x1_txp),
    
        .pcie_perstn         (pcie_perstn),
        .pcie_refclk_clk_n   (pcie_refclk_clk_n),
        .pcie_refclk_clk_p   (pcie_refclk_clk_p),
    
        .qsfp0_156mhz_clk_n  (qsfp0_156mhz_clk_n),
        .qsfp0_156mhz_clk_p  (qsfp0_156mhz_clk_p),
        .qsfp0_1x_grx_n      (qsfp0_1x_grx_n),
        .qsfp0_1x_grx_p      (qsfp0_1x_grx_p),
        .qsfp0_1x_gtx_n      (qsfp0_1x_gtx_n),
        .qsfp0_1x_gtx_p      (qsfp0_1x_gtx_p),
    
        .refclk_300mhz_clk_n (refclk_300mhz_clk_n),
        .refclk_300mhz_clk_p (refclk_300mhz_clk_p)
    );



endmodule

`default_nettype wire