`ifndef PREPROC_REPEAT_H
`define PREPROC_REPEAT_H

/*

This file includes macros which allow for the expansion of repeating
constructs within Verilog and SystemVerilog code. This is based on 
similar methodologies to those used with the C and C++ preprocessor,
namely those features implemented in the BOOST library. The macro as
written supports repeating up to 128 instances, though this file can
be extended to support larger repeating constructs.

Author: Daniel Rozhko, PhD Candidate University of Toronto

*/


`define PP_REPEAT_0(m,d)
`define PP_REPEAT_1(m,d) `m(0,d)
`define PP_REPEAT_2(m,d) `PP_REPEAT_1(m,d) `m(1,d)
`define PP_REPEAT_3(m,d) `PP_REPEAT_2(m,d) `m(2,d)
`define PP_REPEAT_4(m,d) `PP_REPEAT_3(m,d) `m(3,d)
`define PP_REPEAT_5(m,d) `PP_REPEAT_4(m,d) `m(4,d)
`define PP_REPEAT_6(m,d) `PP_REPEAT_5(m,d) `m(5,d)
`define PP_REPEAT_7(m,d) `PP_REPEAT_6(m,d) `m(6,d)
`define PP_REPEAT_8(m,d) `PP_REPEAT_7(m,d) `m(7,d)
`define PP_REPEAT_9(m,d) `PP_REPEAT_8(m,d) `m(8,d)
`define PP_REPEAT_10(m,d) `PP_REPEAT_9(m,d) `m(9,d)
`define PP_REPEAT_11(m,d) `PP_REPEAT_10(m,d) `m(10,d)
`define PP_REPEAT_12(m,d) `PP_REPEAT_11(m,d) `m(11,d)
`define PP_REPEAT_13(m,d) `PP_REPEAT_12(m,d) `m(12,d)
`define PP_REPEAT_14(m,d) `PP_REPEAT_13(m,d) `m(13,d)
`define PP_REPEAT_15(m,d) `PP_REPEAT_14(m,d) `m(14,d)
`define PP_REPEAT_16(m,d) `PP_REPEAT_15(m,d) `m(15,d)
`define PP_REPEAT_17(m,d) `PP_REPEAT_16(m,d) `m(16,d)
`define PP_REPEAT_18(m,d) `PP_REPEAT_17(m,d) `m(17,d)
`define PP_REPEAT_19(m,d) `PP_REPEAT_18(m,d) `m(18,d)
`define PP_REPEAT_20(m,d) `PP_REPEAT_19(m,d) `m(19,d)
`define PP_REPEAT_21(m,d) `PP_REPEAT_20(m,d) `m(20,d)
`define PP_REPEAT_22(m,d) `PP_REPEAT_21(m,d) `m(21,d)
`define PP_REPEAT_23(m,d) `PP_REPEAT_22(m,d) `m(22,d)
`define PP_REPEAT_24(m,d) `PP_REPEAT_23(m,d) `m(23,d)
`define PP_REPEAT_25(m,d) `PP_REPEAT_24(m,d) `m(24,d)
`define PP_REPEAT_26(m,d) `PP_REPEAT_25(m,d) `m(25,d)
`define PP_REPEAT_27(m,d) `PP_REPEAT_26(m,d) `m(26,d)
`define PP_REPEAT_28(m,d) `PP_REPEAT_27(m,d) `m(27,d)
`define PP_REPEAT_29(m,d) `PP_REPEAT_28(m,d) `m(28,d)
`define PP_REPEAT_30(m,d) `PP_REPEAT_29(m,d) `m(29,d)
`define PP_REPEAT_31(m,d) `PP_REPEAT_30(m,d) `m(30,d)
`define PP_REPEAT_32(m,d) `PP_REPEAT_31(m,d) `m(31,d)
`define PP_REPEAT_33(m,d) `PP_REPEAT_32(m,d) `m(32,d)
`define PP_REPEAT_34(m,d) `PP_REPEAT_33(m,d) `m(33,d)
`define PP_REPEAT_35(m,d) `PP_REPEAT_34(m,d) `m(34,d)
`define PP_REPEAT_36(m,d) `PP_REPEAT_35(m,d) `m(35,d)
`define PP_REPEAT_37(m,d) `PP_REPEAT_36(m,d) `m(36,d)
`define PP_REPEAT_38(m,d) `PP_REPEAT_37(m,d) `m(37,d)
`define PP_REPEAT_39(m,d) `PP_REPEAT_38(m,d) `m(38,d)
`define PP_REPEAT_40(m,d) `PP_REPEAT_39(m,d) `m(39,d)
`define PP_REPEAT_41(m,d) `PP_REPEAT_40(m,d) `m(40,d)
`define PP_REPEAT_42(m,d) `PP_REPEAT_41(m,d) `m(41,d)
`define PP_REPEAT_43(m,d) `PP_REPEAT_42(m,d) `m(42,d)
`define PP_REPEAT_44(m,d) `PP_REPEAT_43(m,d) `m(43,d)
`define PP_REPEAT_45(m,d) `PP_REPEAT_44(m,d) `m(44,d)
`define PP_REPEAT_46(m,d) `PP_REPEAT_45(m,d) `m(45,d)
`define PP_REPEAT_47(m,d) `PP_REPEAT_46(m,d) `m(46,d)
`define PP_REPEAT_48(m,d) `PP_REPEAT_47(m,d) `m(47,d)
`define PP_REPEAT_49(m,d) `PP_REPEAT_48(m,d) `m(48,d)
`define PP_REPEAT_50(m,d) `PP_REPEAT_49(m,d) `m(49,d)
`define PP_REPEAT_51(m,d) `PP_REPEAT_50(m,d) `m(50,d)
`define PP_REPEAT_52(m,d) `PP_REPEAT_51(m,d) `m(51,d)
`define PP_REPEAT_53(m,d) `PP_REPEAT_52(m,d) `m(52,d)
`define PP_REPEAT_54(m,d) `PP_REPEAT_53(m,d) `m(53,d)
`define PP_REPEAT_55(m,d) `PP_REPEAT_54(m,d) `m(54,d)
`define PP_REPEAT_56(m,d) `PP_REPEAT_55(m,d) `m(55,d)
`define PP_REPEAT_57(m,d) `PP_REPEAT_56(m,d) `m(56,d)
`define PP_REPEAT_58(m,d) `PP_REPEAT_57(m,d) `m(57,d)
`define PP_REPEAT_59(m,d) `PP_REPEAT_58(m,d) `m(58,d)
`define PP_REPEAT_60(m,d) `PP_REPEAT_59(m,d) `m(59,d)
`define PP_REPEAT_61(m,d) `PP_REPEAT_60(m,d) `m(60,d)
`define PP_REPEAT_62(m,d) `PP_REPEAT_61(m,d) `m(61,d)
`define PP_REPEAT_63(m,d) `PP_REPEAT_62(m,d) `m(62,d)
`define PP_REPEAT_64(m,d) `PP_REPEAT_63(m,d) `m(63,d)
`define PP_REPEAT_65(m,d) `PP_REPEAT_64(m,d) `m(64,d)
`define PP_REPEAT_66(m,d) `PP_REPEAT_65(m,d) `m(65,d)
`define PP_REPEAT_67(m,d) `PP_REPEAT_66(m,d) `m(66,d)
`define PP_REPEAT_68(m,d) `PP_REPEAT_67(m,d) `m(67,d)
`define PP_REPEAT_69(m,d) `PP_REPEAT_68(m,d) `m(68,d)
`define PP_REPEAT_70(m,d) `PP_REPEAT_69(m,d) `m(69,d)
`define PP_REPEAT_71(m,d) `PP_REPEAT_70(m,d) `m(70,d)
`define PP_REPEAT_72(m,d) `PP_REPEAT_71(m,d) `m(71,d)
`define PP_REPEAT_73(m,d) `PP_REPEAT_72(m,d) `m(72,d)
`define PP_REPEAT_74(m,d) `PP_REPEAT_73(m,d) `m(73,d)
`define PP_REPEAT_75(m,d) `PP_REPEAT_74(m,d) `m(74,d)
`define PP_REPEAT_76(m,d) `PP_REPEAT_75(m,d) `m(75,d)
`define PP_REPEAT_77(m,d) `PP_REPEAT_76(m,d) `m(76,d)
`define PP_REPEAT_78(m,d) `PP_REPEAT_77(m,d) `m(77,d)
`define PP_REPEAT_79(m,d) `PP_REPEAT_78(m,d) `m(78,d)
`define PP_REPEAT_80(m,d) `PP_REPEAT_79(m,d) `m(79,d)
`define PP_REPEAT_81(m,d) `PP_REPEAT_80(m,d) `m(80,d)
`define PP_REPEAT_82(m,d) `PP_REPEAT_81(m,d) `m(81,d)
`define PP_REPEAT_83(m,d) `PP_REPEAT_82(m,d) `m(82,d)
`define PP_REPEAT_84(m,d) `PP_REPEAT_83(m,d) `m(83,d)
`define PP_REPEAT_85(m,d) `PP_REPEAT_84(m,d) `m(84,d)
`define PP_REPEAT_86(m,d) `PP_REPEAT_85(m,d) `m(85,d)
`define PP_REPEAT_87(m,d) `PP_REPEAT_86(m,d) `m(86,d)
`define PP_REPEAT_88(m,d) `PP_REPEAT_87(m,d) `m(87,d)
`define PP_REPEAT_89(m,d) `PP_REPEAT_88(m,d) `m(88,d)
`define PP_REPEAT_90(m,d) `PP_REPEAT_89(m,d) `m(89,d)
`define PP_REPEAT_91(m,d) `PP_REPEAT_90(m,d) `m(90,d)
`define PP_REPEAT_92(m,d) `PP_REPEAT_91(m,d) `m(91,d)
`define PP_REPEAT_93(m,d) `PP_REPEAT_92(m,d) `m(92,d)
`define PP_REPEAT_94(m,d) `PP_REPEAT_93(m,d) `m(93,d)
`define PP_REPEAT_95(m,d) `PP_REPEAT_94(m,d) `m(94,d)
`define PP_REPEAT_96(m,d) `PP_REPEAT_95(m,d) `m(95,d)
`define PP_REPEAT_97(m,d) `PP_REPEAT_96(m,d) `m(96,d)
`define PP_REPEAT_98(m,d) `PP_REPEAT_97(m,d) `m(97,d)
`define PP_REPEAT_99(m,d) `PP_REPEAT_98(m,d) `m(98,d)
`define PP_REPEAT_100(m,d) `PP_REPEAT_99(m,d) `m(99,d)
`define PP_REPEAT_101(m,d) `PP_REPEAT_100(m,d) `m(100,d)
`define PP_REPEAT_102(m,d) `PP_REPEAT_101(m,d) `m(101,d)
`define PP_REPEAT_103(m,d) `PP_REPEAT_102(m,d) `m(102,d)
`define PP_REPEAT_104(m,d) `PP_REPEAT_103(m,d) `m(103,d)
`define PP_REPEAT_105(m,d) `PP_REPEAT_104(m,d) `m(104,d)
`define PP_REPEAT_106(m,d) `PP_REPEAT_105(m,d) `m(105,d)
`define PP_REPEAT_107(m,d) `PP_REPEAT_106(m,d) `m(106,d)
`define PP_REPEAT_108(m,d) `PP_REPEAT_107(m,d) `m(107,d)
`define PP_REPEAT_109(m,d) `PP_REPEAT_108(m,d) `m(108,d)
`define PP_REPEAT_110(m,d) `PP_REPEAT_109(m,d) `m(109,d)
`define PP_REPEAT_111(m,d) `PP_REPEAT_110(m,d) `m(110,d)
`define PP_REPEAT_112(m,d) `PP_REPEAT_111(m,d) `m(111,d)
`define PP_REPEAT_113(m,d) `PP_REPEAT_112(m,d) `m(112,d)
`define PP_REPEAT_114(m,d) `PP_REPEAT_113(m,d) `m(113,d)
`define PP_REPEAT_115(m,d) `PP_REPEAT_114(m,d) `m(114,d)
`define PP_REPEAT_116(m,d) `PP_REPEAT_115(m,d) `m(115,d)
`define PP_REPEAT_117(m,d) `PP_REPEAT_116(m,d) `m(116,d)
`define PP_REPEAT_118(m,d) `PP_REPEAT_117(m,d) `m(117,d)
`define PP_REPEAT_119(m,d) `PP_REPEAT_118(m,d) `m(118,d)
`define PP_REPEAT_120(m,d) `PP_REPEAT_119(m,d) `m(119,d)
`define PP_REPEAT_121(m,d) `PP_REPEAT_120(m,d) `m(120,d)
`define PP_REPEAT_122(m,d) `PP_REPEAT_121(m,d) `m(121,d)
`define PP_REPEAT_123(m,d) `PP_REPEAT_122(m,d) `m(122,d)
`define PP_REPEAT_124(m,d) `PP_REPEAT_123(m,d) `m(123,d)
`define PP_REPEAT_125(m,d) `PP_REPEAT_124(m,d) `m(124,d)
`define PP_REPEAT_126(m,d) `PP_REPEAT_125(m,d) `m(125,d)
`define PP_REPEAT_127(m,d) `PP_REPEAT_126(m,d) `m(126,d)
`define PP_REPEAT_128(m,d) `PP_REPEAT_127(m,d) `m(127,d)

`define PP_REPEAT_I(c,m,d) `PP_REPEAT_``c(m,d)
`define PP_REPEAT(c,m,d) `PP_REPEAT_I(c,m,d)


`endif