//Top Level signals to be defined here:

//TODO - update this

  input wire pci_express_x1_rxn,
  input wire pci_express_x1_rxp,
  output wire pci_express_x1_txn,
  output wire pci_express_x1_txp,
  input wire pcie_perstn,
  input wire pcie_refclk_clk_n,
  input wire pcie_refclk_clk_p,
  
  input wire qsfp0_156mhz_clk_n,
  input wire qsfp0_156mhz_clk_p,
  input wire qsfp0_1x_grx_n,
  input wire qsfp0_1x_grx_p,
  output wire qsfp0_1x_gtx_n,
  output wire qsfp0_1x_gtx_p,
  input wire refclk_300mhz_clk_n,
  input wire refclk_300mhz_clk_p