`timescale 1ns / 1ps
`default_nettype none

/*
Shell Wrapper for physical layer interfaces (to be implemented per platform)

Author: Daniel Rozhko, PhD Candidate University of Toronto

Description:
   This module wraps all of the physcial layer interfaces needed by the
   shell, which includes a network interface (TX and RX) and some control 
   interface (e.g. PCIe).

Parameters:
   NET_AXIS_BUS_WIDTH - the data width of the axi-streams (must be multiple of 8)
   NET_MAX_PACKET_LENGTH - the maximum network packet length to support (for forced tlast)

Ports:
   axis_tx_s_* - the input axi stream for the tx direction, to phy
   axis_rx_m_* - the output axi stream for the rx direction, from phy
   axis_aclk - clock to which all of the network signals are synchronous (generated by physical layer)
   axis_aresetn - active-low reset corresponding to above clock (generated by physical layer)

   top_ctrl_* - the AXI-Lite control interface for the top-level control (e.g. PCIe)
   top_mem_* - the AXI4 memory-access interface for the top-level (e.g. PCIe)
   top_aclk - clock to which the control signal is synchronous (generated by physical layer)
   top_aresetn - active-low reset corresponding to above clock (generated by physical layer)

Notes:
   - Various portions of the hdl below require the manual addition of vendor
   specific cores for clock crossing and AXI switching/crossbar. Search for 
   [VENDOR SPECIFIC] for all places where such cores are required
   - all platform specific ports need to be added to the file for each platform
   implementation
*/


module phy_shell
#(
    //Network AXI Stream Params (as seen by application regions)
    parameter NET_AXIS_BUS_WIDTH = 64,

    //Network Packet Params
    parameter NET_MAX_PACKET_LENGTH = 1522



    //AXI-Lite Interface Params
    //parameter CTRL_AXI_DATA_WIDTH = 32, //Fixed to 32 for now, 64-bit not supported by some cores
)
(
    //Egress Output AXI stream (TX packets to Phy)
    input wire [NET_AXIS_BUS_WIDTH-1:0]          axis_tx_s_tdata,
    input wire [(NET_AXIS_BUS_WIDTH/8)-1:0]      axis_tx_s_tkeep,
    input wire                                   axis_tx_s_tlast,
    input wire                                   axis_tx_s_tvalid,
    output wire                                  axis_tx_s_tready,

    //Ingress Input AXI stream (RX packets from Phy)
    output wire [NET_AXIS_BUS_WIDTH-1:0]         axis_rx_m_tdata,
    output wire [(NET_AXIS_BUS_WIDTH/8)-1:0]     axis_rx_m_tkeep,
    output wire                                  axis_rx_m_tlast,
    output wire                                  axis_rx_m_tvalid,
    input wire                                   axis_rx_m_tready,

    //Network Clocking
    output wire  axis_aclk,
    output wire  axis_aresetn,
    


    //The AXI-Lite Control Interface (from control, e.g. PCIe)
    //Write Address Channel  
    output wire  [31:0]                        top_ctrl_awaddr,
    output wire                                top_ctrl_awvalid,
    input wire                                 top_ctrl_awready,
    //Write Data Channel
    output wire  [31:0]                        top_ctrl_wdata,
    output wire  [3:0]                         top_ctrl_wstrb,
    output wire                                top_ctrl_wvalid,
    input wire                                 top_ctrl_wready,
    //Write Response Channel
    input wire [1:0]                           top_ctrl_bresp,
    input wire                                 top_ctrl_bvalid,
    output wire                                top_ctrl_bready,
    //Read Address Channel 
    output wire  [31:0]                        top_ctrl_araddr,
    output wire                                top_ctrl_arvalid,
    input wire                                 top_ctrl_arready,
    //Read Data Response Channel
    input wire [31:0]                          top_ctrl_rdata,
    input wire [1:0]                           top_ctrl_rresp,
    input wire                                 top_ctrl_rvalid,
    output wire                                top_ctrl_rready,

    //Ctrl Clocking
    output wire  top_aclk,
    output wire  top_aresetn,
    
    //Physical layer ports (from include file)
    `include "phy_signals.svh"
);

    //--------------------------------------------------------//
    //   PHY for network access                               //
    //--------------------------------------------------------//

    //[VENDOR SPECIFIC]
    //Insert the vencor specific network PHY (e.g. 10G Ethernet Controller)
    //   - Input interface for tx is axis_tx_s_*, sync to axis_aclk
    //   - Output interafce for tx is the pins added above (platform specific)
    //   - Input interface for rx is the pins added above (platform specific)
    //   - Output interface for rx is axis_rx_m_*, sync to axis_aclk
    //       - note, no tready (no back pressure)
    //   - The clock signals axis_aclk and axis_aresetn should be driven here 




    //--------------------------------------------------------//
    //   PHY for control access (e.g. PCIe)                   //
    //--------------------------------------------------------//

    //[VENDOR SPECIFIC]
    //Insert the vencor specific control PHY (e.g. PCIe XDMA)
    //   - Input interafce is the pins added above (platform specific)
    //   - Output interface for control is top_ctrl_*, sync to top_aclk
    //   - The clock signals top_aclk and top_aresetn should be driven here 




endmodule

`default_nettype wire