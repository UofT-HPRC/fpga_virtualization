`timescale 1ns / 1ps
`default_nettype none


//Number of masters
`define NUM_MASTERS 4
`define INC_M1
`define INC_M2
`define INC_M3
`define INC_M4
//`define INC_M5
//`define INC_M6
//`define INC_M7
//`define INC_M8

//The memory prtocol checker/corrector
module mem_bw_throttler_multi_wrapper
#(
    //AXI4 Interface Params
    parameter AXI_ID_WIDTH = 4,
    parameter AXI_ADDR_WIDTH = 32,
    parameter AXI_DATA_WIDTH = 128,
    parameter AXI_AX_USER_WIDTH = 1,
    
    //Token counter params
    parameter TOKEN_COUNT_INT_WIDTH = 16,
    parameter TOKEN_COUNT_FRAC_WIDTH = 8,
    localparam BW_THROT_BITS_PER_MAST = (TOKEN_COUNT_INT_WIDTH + TOKEN_COUNT_FRAC_WIDTH + 1) * 2,
    localparam BW_THROT_REG_WIDTH =  BW_THROT_BITS_PER_MAST * `NUM_MASTERS,

    //Timeout limits
    parameter WTIMEOUT_CYCLES = 15,
    parameter BTIMEOUT_CYCLES = 15,
    parameter RTIMEOUT_CYCLES = 15,
    parameter OUTSTANDING_WREQ = 8,
    parameter OUTSTANDING_RREQ = 8,

    //Retiming for adders
    parameter AW_RETIMING_STAGES = 0,
    parameter AR_RETIMING_STAGES = 0,

    //Features to Implement
    parameter ALLOW_OVERRIDE = 1,
    parameter INCLUDE_BACKPRESSURE = 0
)
(

`ifdef INC_M1

    //AXI4 slave connection (input of requests)
    //Write Address Channel
    input wire [AXI_ID_WIDTH-1:0]           in1_awid,
    input wire [AXI_ADDR_WIDTH-1:0]         in1_awaddr,
    input wire [7:0]                        in1_awlen,
    input wire [2:0]                        in1_awsize,
    input wire [1:0]                        in1_awburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in1_awuser,
    input wire                              in1_awvalid,
    output wire                             in1_awready,
    //Write Data Channel
    input wire [AXI_DATA_WIDTH-1:0]         in1_wdata,
    input wire [(AXI_DATA_WIDTH/8)-1:0]     in1_wstrb,
    input wire                              in1_wlast,
    input wire                              in1_wvalid,
    output wire                             in1_wready,
    //Write Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in1_bid,
    output wire [1:0]                       in1_bresp,
    output wire                             in1_bvalid,
    input wire                              in1_bready,
    //Read Address Channel     
    input wire [AXI_ID_WIDTH-1:0]           in1_arid,
    input wire [AXI_ADDR_WIDTH-1:0]         in1_araddr,
    input wire [7:0]                        in1_arlen,
    input wire [2:0]                        in1_arsize,
    input wire [1:0]                        in1_arburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in1_aruser,
    input wire                              in1_arvalid,
    output wire                             in1_arready,
    //Read Data Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in1_rid,
    output wire [AXI_DATA_WIDTH-1:0]        in1_rdata,
    output wire [1:0]                       in1_rresp,
    output wire                             in1_rlast,
    output wire                             in1_rvalid,
    input wire                              in1_rready,

    //AXI4 master connection (output of requests)
    //Write Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out1_awid,
    output wire [AXI_ADDR_WIDTH-1:0]        out1_awaddr,
    output wire [7:0]                       out1_awlen,
    output wire [2:0]                       out1_awsize,
    output wire [1:0]                       out1_awburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out1_awuser,
    output wire                             out1_awvalid,
    input wire                              out1_awready,
    //Write Data Channel
    output wire [AXI_DATA_WIDTH-1:0]        out1_wdata,
    output wire [(AXI_DATA_WIDTH/8)-1:0]    out1_wstrb,
    output wire                             out1_wlast,
    output wire                             out1_wvalid,
    input wire                              out1_wready,
    //Write Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out1_bid,
    input wire [1:0]                        out1_bresp,
    input wire                              out1_bvalid,
    output wire                             out1_bready,
    //Read Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out1_arid,
    output wire [AXI_ADDR_WIDTH-1:0]        out1_araddr,
    output wire [7:0]                       out1_arlen,
    output wire [2:0]                       out1_arsize,
    output wire [1:0]                       out1_arburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out1_aruser,
    output wire                             out1_arvalid,
    input wire                              out1_arready,
    //Read Data Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out1_rid,
    input wire [AXI_DATA_WIDTH-1:0]         out1_rdata,
    input wire [1:0]                        out1_rresp,
    input wire                              out1_rlast,
    input wire                              out1_rvalid,
    output wire                             out1_rready,

`endif

`ifdef INC_M2

    //AXI4 slave connection (input of requests)
    //Write Address Channel
    input wire [AXI_ID_WIDTH-1:0]           in2_awid,
    input wire [AXI_ADDR_WIDTH-1:0]         in2_awaddr,
    input wire [7:0]                        in2_awlen,
    input wire [2:0]                        in2_awsize,
    input wire [1:0]                        in2_awburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in2_awuser,
    input wire                              in2_awvalid,
    output wire                             in2_awready,
    //Write Data Channel
    input wire [AXI_DATA_WIDTH-1:0]         in2_wdata,
    input wire [(AXI_DATA_WIDTH/8)-1:0]     in2_wstrb,
    input wire                              in2_wlast,
    input wire                              in2_wvalid,
    output wire                             in2_wready,
    //Write Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in2_bid,
    output wire [1:0]                       in2_bresp,
    output wire                             in2_bvalid,
    input wire                              in2_bready,
    //Read Address Channel     
    input wire [AXI_ID_WIDTH-1:0]           in2_arid,
    input wire [AXI_ADDR_WIDTH-1:0]         in2_araddr,
    input wire [7:0]                        in2_arlen,
    input wire [2:0]                        in2_arsize,
    input wire [1:0]                        in2_arburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in2_aruser,
    input wire                              in2_arvalid,
    output wire                             in2_arready,
    //Read Data Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in2_rid,
    output wire [AXI_DATA_WIDTH-1:0]        in2_rdata,
    output wire [1:0]                       in2_rresp,
    output wire                             in2_rlast,
    output wire                             in2_rvalid,
    input wire                              in2_rready,

    //AXI4 master connection (output of requests)
    //Write Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out2_awid,
    output wire [AXI_ADDR_WIDTH-1:0]        out2_awaddr,
    output wire [7:0]                       out2_awlen,
    output wire [2:0]                       out2_awsize,
    output wire [1:0]                       out2_awburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out2_awuser,
    output wire                             out2_awvalid,
    input wire                              out2_awready,
    //Write Data Channel
    output wire [AXI_DATA_WIDTH-1:0]        out2_wdata,
    output wire [(AXI_DATA_WIDTH/8)-1:0]    out2_wstrb,
    output wire                             out2_wlast,
    output wire                             out2_wvalid,
    input wire                              out2_wready,
    //Write Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out2_bid,
    input wire [1:0]                        out2_bresp,
    input wire                              out2_bvalid,
    output wire                             out2_bready,
    //Read Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out2_arid,
    output wire [AXI_ADDR_WIDTH-1:0]        out2_araddr,
    output wire [7:0]                       out2_arlen,
    output wire [2:0]                       out2_arsize,
    output wire [1:0]                       out2_arburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out2_aruser,
    output wire                             out2_arvalid,
    input wire                              out2_arready,
    //Read Data Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out2_rid,
    input wire [AXI_DATA_WIDTH-1:0]         out2_rdata,
    input wire [1:0]                        out2_rresp,
    input wire                              out2_rlast,
    input wire                              out2_rvalid,
    output wire                             out2_rready,

`endif

`ifdef INC_M3

    //AXI4 slave connection (input of requests)
    //Write Address Channel
    input wire [AXI_ID_WIDTH-1:0]           in3_awid,
    input wire [AXI_ADDR_WIDTH-1:0]         in3_awaddr,
    input wire [7:0]                        in3_awlen,
    input wire [2:0]                        in3_awsize,
    input wire [1:0]                        in3_awburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in3_awuser,
    input wire                              in3_awvalid,
    output wire                             in3_awready,
    //Write Data Channel
    input wire [AXI_DATA_WIDTH-1:0]         in3_wdata,
    input wire [(AXI_DATA_WIDTH/8)-1:0]     in3_wstrb,
    input wire                              in3_wlast,
    input wire                              in3_wvalid,
    output wire                             in3_wready,
    //Write Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in3_bid,
    output wire [1:0]                       in3_bresp,
    output wire                             in3_bvalid,
    input wire                              in3_bready,
    //Read Address Channel     
    input wire [AXI_ID_WIDTH-1:0]           in3_arid,
    input wire [AXI_ADDR_WIDTH-1:0]         in3_araddr,
    input wire [7:0]                        in3_arlen,
    input wire [2:0]                        in3_arsize,
    input wire [1:0]                        in3_arburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in3_aruser,
    input wire                              in3_arvalid,
    output wire                             in3_arready,
    //Read Data Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in3_rid,
    output wire [AXI_DATA_WIDTH-1:0]        in3_rdata,
    output wire [1:0]                       in3_rresp,
    output wire                             in3_rlast,
    output wire                             in3_rvalid,
    input wire                              in3_rready,

    //AXI4 master connection (output of requests)
    //Write Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out3_awid,
    output wire [AXI_ADDR_WIDTH-1:0]        out3_awaddr,
    output wire [7:0]                       out3_awlen,
    output wire [2:0]                       out3_awsize,
    output wire [1:0]                       out3_awburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out3_awuser,
    output wire                             out3_awvalid,
    input wire                              out3_awready,
    //Write Data Channel
    output wire [AXI_DATA_WIDTH-1:0]        out3_wdata,
    output wire [(AXI_DATA_WIDTH/8)-1:0]    out3_wstrb,
    output wire                             out3_wlast,
    output wire                             out3_wvalid,
    input wire                              out3_wready,
    //Write Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out3_bid,
    input wire [1:0]                        out3_bresp,
    input wire                              out3_bvalid,
    output wire                             out3_bready,
    //Read Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out3_arid,
    output wire [AXI_ADDR_WIDTH-1:0]        out3_araddr,
    output wire [7:0]                       out3_arlen,
    output wire [2:0]                       out3_arsize,
    output wire [1:0]                       out3_arburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out3_aruser,
    output wire                             out3_arvalid,
    input wire                              out3_arready,
    //Read Data Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out3_rid,
    input wire [AXI_DATA_WIDTH-1:0]         out3_rdata,
    input wire [1:0]                        out3_rresp,
    input wire                              out3_rlast,
    input wire                              out3_rvalid,
    output wire                             out3_rready,

`endif

`ifdef INC_M4

    //AXI4 slave connection (input of requests)
    //Write Address Channel
    input wire [AXI_ID_WIDTH-1:0]           in4_awid,
    input wire [AXI_ADDR_WIDTH-1:0]         in4_awaddr,
    input wire [7:0]                        in4_awlen,
    input wire [2:0]                        in4_awsize,
    input wire [1:0]                        in4_awburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in4_awuser,
    input wire                              in4_awvalid,
    output wire                             in4_awready,
    //Write Data Channel
    input wire [AXI_DATA_WIDTH-1:0]         in4_wdata,
    input wire [(AXI_DATA_WIDTH/8)-1:0]     in4_wstrb,
    input wire                              in4_wlast,
    input wire                              in4_wvalid,
    output wire                             in4_wready,
    //Write Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in4_bid,
    output wire [1:0]                       in4_bresp,
    output wire                             in4_bvalid,
    input wire                              in4_bready,
    //Read Address Channel     
    input wire [AXI_ID_WIDTH-1:0]           in4_arid,
    input wire [AXI_ADDR_WIDTH-1:0]         in4_araddr,
    input wire [7:0]                        in4_arlen,
    input wire [2:0]                        in4_arsize,
    input wire [1:0]                        in4_arburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in4_aruser,
    input wire                              in4_arvalid,
    output wire                             in4_arready,
    //Read Data Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in4_rid,
    output wire [AXI_DATA_WIDTH-1:0]        in4_rdata,
    output wire [1:0]                       in4_rresp,
    output wire                             in4_rlast,
    output wire                             in4_rvalid,
    input wire                              in4_rready,

    //AXI4 master connection (output of requests)
    //Write Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out4_awid,
    output wire [AXI_ADDR_WIDTH-1:0]        out4_awaddr,
    output wire [7:0]                       out4_awlen,
    output wire [2:0]                       out4_awsize,
    output wire [1:0]                       out4_awburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out4_awuser,
    output wire                             out4_awvalid,
    input wire                              out4_awready,
    //Write Data Channel
    output wire [AXI_DATA_WIDTH-1:0]        out4_wdata,
    output wire [(AXI_DATA_WIDTH/8)-1:0]    out4_wstrb,
    output wire                             out4_wlast,
    output wire                             out4_wvalid,
    input wire                              out4_wready,
    //Write Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out4_bid,
    input wire [1:0]                        out4_bresp,
    input wire                              out4_bvalid,
    output wire                             out4_bready,
    //Read Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out4_arid,
    output wire [AXI_ADDR_WIDTH-1:0]        out4_araddr,
    output wire [7:0]                       out4_arlen,
    output wire [2:0]                       out4_arsize,
    output wire [1:0]                       out4_arburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out4_aruser,
    output wire                             out4_arvalid,
    input wire                              out4_arready,
    //Read Data Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out4_rid,
    input wire [AXI_DATA_WIDTH-1:0]         out4_rdata,
    input wire [1:0]                        out4_rresp,
    input wire                              out4_rlast,
    input wire                              out4_rvalid,
    output wire                             out4_rready,

`endif

`ifdef INC_M5

    //AXI4 slave connection (input of requests)
    //Write Address Channel
    input wire [AXI_ID_WIDTH-1:0]           in5_awid,
    input wire [AXI_ADDR_WIDTH-1:0]         in5_awaddr,
    input wire [7:0]                        in5_awlen,
    input wire [2:0]                        in5_awsize,
    input wire [1:0]                        in5_awburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in5_awuser,
    input wire                              in5_awvalid,
    output wire                             in5_awready,
    //Write Data Channel
    input wire [AXI_DATA_WIDTH-1:0]         in5_wdata,
    input wire [(AXI_DATA_WIDTH/8)-1:0]     in5_wstrb,
    input wire                              in5_wlast,
    input wire                              in5_wvalid,
    output wire                             in5_wready,
    //Write Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in5_bid,
    output wire [1:0]                       in5_bresp,
    output wire                             in5_bvalid,
    input wire                              in5_bready,
    //Read Address Channel     
    input wire [AXI_ID_WIDTH-1:0]           in5_arid,
    input wire [AXI_ADDR_WIDTH-1:0]         in5_araddr,
    input wire [7:0]                        in5_arlen,
    input wire [2:0]                        in5_arsize,
    input wire [1:0]                        in5_arburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in5_aruser,
    input wire                              in5_arvalid,
    output wire                             in5_arready,
    //Read Data Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in5_rid,
    output wire [AXI_DATA_WIDTH-1:0]        in5_rdata,
    output wire [1:0]                       in5_rresp,
    output wire                             in5_rlast,
    output wire                             in5_rvalid,
    input wire                              in5_rready,

    //AXI4 master connection (output of requests)
    //Write Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out5_awid,
    output wire [AXI_ADDR_WIDTH-1:0]        out5_awaddr,
    output wire [7:0]                       out5_awlen,
    output wire [2:0]                       out5_awsize,
    output wire [1:0]                       out5_awburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out5_awuser,
    output wire                             out5_awvalid,
    input wire                              out5_awready,
    //Write Data Channel
    output wire [AXI_DATA_WIDTH-1:0]        out5_wdata,
    output wire [(AXI_DATA_WIDTH/8)-1:0]    out5_wstrb,
    output wire                             out5_wlast,
    output wire                             out5_wvalid,
    input wire                              out5_wready,
    //Write Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out5_bid,
    input wire [1:0]                        out5_bresp,
    input wire                              out5_bvalid,
    output wire                             out5_bready,
    //Read Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out5_arid,
    output wire [AXI_ADDR_WIDTH-1:0]        out5_araddr,
    output wire [7:0]                       out5_arlen,
    output wire [2:0]                       out5_arsize,
    output wire [1:0]                       out5_arburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out5_aruser,
    output wire                             out5_arvalid,
    input wire                              out5_arready,
    //Read Data Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out5_rid,
    input wire [AXI_DATA_WIDTH-1:0]         out5_rdata,
    input wire [1:0]                        out5_rresp,
    input wire                              out5_rlast,
    input wire                              out5_rvalid,
    output wire                             out5_rready,

`endif

`ifdef INC_M6

    //AXI4 slave connection (input of requests)
    //Write Address Channel
    input wire [AXI_ID_WIDTH-1:0]           in6_awid,
    input wire [AXI_ADDR_WIDTH-1:0]         in6_awaddr,
    input wire [7:0]                        in6_awlen,
    input wire [2:0]                        in6_awsize,
    input wire [1:0]                        in6_awburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in6_awuser,
    input wire                              in6_awvalid,
    output wire                             in6_awready,
    //Write Data Channel
    input wire [AXI_DATA_WIDTH-1:0]         in6_wdata,
    input wire [(AXI_DATA_WIDTH/8)-1:0]     in6_wstrb,
    input wire                              in6_wlast,
    input wire                              in6_wvalid,
    output wire                             in6_wready,
    //Write Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in6_bid,
    output wire [1:0]                       in6_bresp,
    output wire                             in6_bvalid,
    input wire                              in6_bready,
    //Read Address Channel     
    input wire [AXI_ID_WIDTH-1:0]           in6_arid,
    input wire [AXI_ADDR_WIDTH-1:0]         in6_araddr,
    input wire [7:0]                        in6_arlen,
    input wire [2:0]                        in6_arsize,
    input wire [1:0]                        in6_arburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in6_aruser,
    input wire                              in6_arvalid,
    output wire                             in6_arready,
    //Read Data Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in6_rid,
    output wire [AXI_DATA_WIDTH-1:0]        in6_rdata,
    output wire [1:0]                       in6_rresp,
    output wire                             in6_rlast,
    output wire                             in6_rvalid,
    input wire                              in6_rready,

    //AXI4 master connection (output of requests)
    //Write Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out6_awid,
    output wire [AXI_ADDR_WIDTH-1:0]        out6_awaddr,
    output wire [7:0]                       out6_awlen,
    output wire [2:0]                       out6_awsize,
    output wire [1:0]                       out6_awburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out6_awuser,
    output wire                             out6_awvalid,
    input wire                              out6_awready,
    //Write Data Channel
    output wire [AXI_DATA_WIDTH-1:0]        out6_wdata,
    output wire [(AXI_DATA_WIDTH/8)-1:0]    out6_wstrb,
    output wire                             out6_wlast,
    output wire                             out6_wvalid,
    input wire                              out6_wready,
    //Write Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out6_bid,
    input wire [1:0]                        out6_bresp,
    input wire                              out6_bvalid,
    output wire                             out6_bready,
    //Read Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out6_arid,
    output wire [AXI_ADDR_WIDTH-1:0]        out6_araddr,
    output wire [7:0]                       out6_arlen,
    output wire [2:0]                       out6_arsize,
    output wire [1:0]                       out6_arburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out6_aruser,
    output wire                             out6_arvalid,
    input wire                              out6_arready,
    //Read Data Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out6_rid,
    input wire [AXI_DATA_WIDTH-1:0]         out6_rdata,
    input wire [1:0]                        out6_rresp,
    input wire                              out6_rlast,
    input wire                              out6_rvalid,
    output wire                             out6_rready,

`endif

`ifdef INC_M7

    //AXI4 slave connection (input of requests)
    //Write Address Channel
    input wire [AXI_ID_WIDTH-1:0]           in7_awid,
    input wire [AXI_ADDR_WIDTH-1:0]         in7_awaddr,
    input wire [7:0]                        in7_awlen,
    input wire [2:0]                        in7_awsize,
    input wire [1:0]                        in7_awburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in7_awuser,
    input wire                              in7_awvalid,
    output wire                             in7_awready,
    //Write Data Channel
    input wire [AXI_DATA_WIDTH-1:0]         in7_wdata,
    input wire [(AXI_DATA_WIDTH/8)-1:0]     in7_wstrb,
    input wire                              in7_wlast,
    input wire                              in7_wvalid,
    output wire                             in7_wready,
    //Write Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in7_bid,
    output wire [1:0]                       in7_bresp,
    output wire                             in7_bvalid,
    input wire                              in7_bready,
    //Read Address Channel     
    input wire [AXI_ID_WIDTH-1:0]           in7_arid,
    input wire [AXI_ADDR_WIDTH-1:0]         in7_araddr,
    input wire [7:0]                        in7_arlen,
    input wire [2:0]                        in7_arsize,
    input wire [1:0]                        in7_arburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in7_aruser,
    input wire                              in7_arvalid,
    output wire                             in7_arready,
    //Read Data Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in7_rid,
    output wire [AXI_DATA_WIDTH-1:0]        in7_rdata,
    output wire [1:0]                       in7_rresp,
    output wire                             in7_rlast,
    output wire                             in7_rvalid,
    input wire                              in7_rready,

    //AXI4 master connection (output of requests)
    //Write Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out7_awid,
    output wire [AXI_ADDR_WIDTH-1:0]        out7_awaddr,
    output wire [7:0]                       out7_awlen,
    output wire [2:0]                       out7_awsize,
    output wire [1:0]                       out7_awburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out7_awuser,
    output wire                             out7_awvalid,
    input wire                              out7_awready,
    //Write Data Channel
    output wire [AXI_DATA_WIDTH-1:0]        out7_wdata,
    output wire [(AXI_DATA_WIDTH/8)-1:0]    out7_wstrb,
    output wire                             out7_wlast,
    output wire                             out7_wvalid,
    input wire                              out7_wready,
    //Write Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out7_bid,
    input wire [1:0]                        out7_bresp,
    input wire                              out7_bvalid,
    output wire                             out7_bready,
    //Read Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out7_arid,
    output wire [AXI_ADDR_WIDTH-1:0]        out7_araddr,
    output wire [7:0]                       out7_arlen,
    output wire [2:0]                       out7_arsize,
    output wire [1:0]                       out7_arburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out7_aruser,
    output wire                             out7_arvalid,
    input wire                              out7_arready,
    //Read Data Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out7_rid,
    input wire [AXI_DATA_WIDTH-1:0]         out7_rdata,
    input wire [1:0]                        out7_rresp,
    input wire                              out7_rlast,
    input wire                              out7_rvalid,
    output wire                             out7_rready,

`endif

`ifdef INC_M8

    //AXI4 slave connection (input of requests)
    //Write Address Channel
    input wire [AXI_ID_WIDTH-1:0]           in8_awid,
    input wire [AXI_ADDR_WIDTH-1:0]         in8_awaddr,
    input wire [7:0]                        in8_awlen,
    input wire [2:0]                        in8_awsize,
    input wire [1:0]                        in8_awburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in8_awuser,
    input wire                              in8_awvalid,
    output wire                             in8_awready,
    //Write Data Channel
    input wire [AXI_DATA_WIDTH-1:0]         in8_wdata,
    input wire [(AXI_DATA_WIDTH/8)-1:0]     in8_wstrb,
    input wire                              in8_wlast,
    input wire                              in8_wvalid,
    output wire                             in8_wready,
    //Write Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in8_bid,
    output wire [1:0]                       in8_bresp,
    output wire                             in8_bvalid,
    input wire                              in8_bready,
    //Read Address Channel     
    input wire [AXI_ID_WIDTH-1:0]           in8_arid,
    input wire [AXI_ADDR_WIDTH-1:0]         in8_araddr,
    input wire [7:0]                        in8_arlen,
    input wire [2:0]                        in8_arsize,
    input wire [1:0]                        in8_arburst,
    input wire [AXI_AX_USER_WIDTH-1:0]      in8_aruser,
    input wire                              in8_arvalid,
    output wire                             in8_arready,
    //Read Data Response Channel
    output wire [AXI_ID_WIDTH-1:0]          in8_rid,
    output wire [AXI_DATA_WIDTH-1:0]        in8_rdata,
    output wire [1:0]                       in8_rresp,
    output wire                             in8_rlast,
    output wire                             in8_rvalid,
    input wire                              in8_rready,

    //AXI4 master connection (output of requests)
    //Write Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out8_awid,
    output wire [AXI_ADDR_WIDTH-1:0]        out8_awaddr,
    output wire [7:0]                       out8_awlen,
    output wire [2:0]                       out8_awsize,
    output wire [1:0]                       out8_awburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out8_awuser,
    output wire                             out8_awvalid,
    input wire                              out8_awready,
    //Write Data Channel
    output wire [AXI_DATA_WIDTH-1:0]        out8_wdata,
    output wire [(AXI_DATA_WIDTH/8)-1:0]    out8_wstrb,
    output wire                             out8_wlast,
    output wire                             out8_wvalid,
    input wire                              out8_wready,
    //Write Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out8_bid,
    input wire [1:0]                        out8_bresp,
    input wire                              out8_bvalid,
    output wire                             out8_bready,
    //Read Address Channel     
    output wire [AXI_ID_WIDTH-1:0]          out8_arid,
    output wire [AXI_ADDR_WIDTH-1:0]        out8_araddr,
    output wire [7:0]                       out8_arlen,
    output wire [2:0]                       out8_arsize,
    output wire [1:0]                       out8_arburst,
    output wire [AXI_AX_USER_WIDTH-1:0]     out8_aruser,
    output wire                             out8_arvalid,
    input wire                              out8_arready,
    //Read Data Response Channel
    input wire [AXI_ID_WIDTH-1:0]           out8_rid,
    input wire [AXI_DATA_WIDTH-1:0]         out8_rdata,
    input wire [1:0]                        out8_rresp,
    input wire                              out8_rlast,
    input wire                              out8_rvalid,
    output wire                             out8_rready,

`endif

    //Packed Register signals
    input wire [((TOKEN_COUNT_INT_WIDTH+TOKEN_COUNT_FRAC_WIDTH+1)*2*`NUM_MASTERS)-1:0]     
                                            bw_throt_regs,

    //Clocking
    input wire  aclk,
    input wire  aresetn
);


    mem_bw_throttler_multi_wrap_sv
    #(
        .AXI_ID_WIDTH           (AXI_ID_WIDTH),
        .AXI_ADDR_WIDTH         (AXI_ADDR_WIDTH),
        .AXI_DATA_WIDTH         (AXI_DATA_WIDTH),
        .AXI_AX_USER_WIDTH      (AXI_AX_USER_WIDTH),
        .TOKEN_COUNT_INT_WIDTH  (TOKEN_COUNT_INT_WIDTH),
        .TOKEN_COUNT_FRAC_WIDTH (TOKEN_COUNT_FRAC_WIDTH),
        .WTIMEOUT_CYCLES        (WTIMEOUT_CYCLES),
        .BTIMEOUT_CYCLES        (BTIMEOUT_CYCLES),
        .RTIMEOUT_CYCLES        (RTIMEOUT_CYCLES),
        .OUTSTANDING_WREQ       (OUTSTANDING_WREQ),
        .OUTSTANDING_RREQ       (OUTSTANDING_RREQ),
        .AW_RETIMING_STAGES     (AW_RETIMING_STAGES),
        .AR_RETIMING_STAGES     (AR_RETIMING_STAGES),
        .ALLOW_OVERRIDE         (ALLOW_OVERRIDE),
        .INCLUDE_BACKPRESSURE   (INCLUDE_BACKPRESSURE)
    )
    thottles 
    (
        
    `ifdef INC_M1

        .in1_awid (in1_awid),
        .in1_awaddr (in1_awaddr),
        .in1_awlen (in1_awlen),
        .in1_awsize (in1_awsize),
        .in1_awburst (in1_awburst),
        .in1_awuser (in1_awuser),
        .in1_awvalid (in1_awvalid),
        .in1_awready (in1_awready),
        .in1_wdata (in1_wdata),
        .in1_wstrb (in1_wstrb),
        .in1_wlast (in1_wlast),
        .in1_wvalid (in1_wvalid),
        .in1_wready (in1_wready),
        .in1_bid (in1_bid),
        .in1_bresp (in1_bresp),
        .in1_bvalid (in1_bvalid),
        .in1_bready (in1_bready),
        .in1_arid (in1_arid),
        .in1_araddr (in1_araddr),
        .in1_arlen (in1_arlen),
        .in1_arsize (in1_arsize),
        .in1_arburst (in1_arburst),
        .in1_aruser (in1_aruser),
        .in1_arvalid (in1_arvalid),
        .in1_arready (in1_arready),
        .in1_rid (in1_rid),
        .in1_rdata (in1_rdata),
        .in1_rresp (in1_rresp),
        .in1_rlast (in1_rlast),
        .in1_rvalid (in1_rvalid),
        .in1_rready (in1_rready),

        .out1_awid (out1_awid),
        .out1_awaddr (out1_awaddr),
        .out1_awlen (out1_awlen),
        .out1_awsize (out1_awsize),
        .out1_awburst (out1_awburst),
        .out1_awuser (out1_awuser),
        .out1_awvalid (out1_awvalid),
        .out1_awready (out1_awready),
        .out1_wdata (out1_wdata),
        .out1_wstrb (out1_wstrb),
        .out1_wlast (out1_wlast),
        .out1_wvalid (out1_wvalid),
        .out1_wready (out1_wready),
        .out1_bid (out1_bid),
        .out1_bresp (out1_bresp),
        .out1_bvalid (out1_bvalid),
        .out1_bready (out1_bready),
        .out1_arid (out1_arid),
        .out1_araddr (out1_araddr),
        .out1_arlen (out1_arlen),
        .out1_arsize (out1_arsize),
        .out1_arburst (out1_arburst),
        .out1_aruser (out1_aruser),
        .out1_arvalid (out1_arvalid),
        .out1_arready (out1_arready),
        .out1_rid (out1_rid),
        .out1_rdata (out1_rdata),
        .out1_rresp (out1_rresp),
        .out1_rlast (out1_rlast),
        .out1_rvalid (out1_rvalid),
        .out1_rready (out1_rready),

    `endif

    `ifdef INC_M2

        .in2_awid (in2_awid),
        .in2_awaddr (in2_awaddr),
        .in2_awlen (in2_awlen),
        .in2_awsize (in2_awsize),
        .in2_awburst (in2_awburst),
        .in2_awuser (in2_awuser),
        .in2_awvalid (in2_awvalid),
        .in2_awready (in2_awready),
        .in2_wdata (in2_wdata),
        .in2_wstrb (in2_wstrb),
        .in2_wlast (in2_wlast),
        .in2_wvalid (in2_wvalid),
        .in2_wready (in2_wready),
        .in2_bid (in2_bid),
        .in2_bresp (in2_bresp),
        .in2_bvalid (in2_bvalid),
        .in2_bready (in2_bready),
        .in2_arid (in2_arid),
        .in2_araddr (in2_araddr),
        .in2_arlen (in2_arlen),
        .in2_arsize (in2_arsize),
        .in2_arburst (in2_arburst),
        .in2_aruser (in2_aruser),
        .in2_arvalid (in2_arvalid),
        .in2_arready (in2_arready),
        .in2_rid (in2_rid),
        .in2_rdata (in2_rdata),
        .in2_rresp (in2_rresp),
        .in2_rlast (in2_rlast),
        .in2_rvalid (in2_rvalid),
        .in2_rready (in2_rready),

        .out2_awid (out2_awid),
        .out2_awaddr (out2_awaddr),
        .out2_awlen (out2_awlen),
        .out2_awsize (out2_awsize),
        .out2_awburst (out2_awburst),
        .out2_awuser (out2_awuser),
        .out2_awvalid (out2_awvalid),
        .out2_awready (out2_awready),
        .out2_wdata (out2_wdata),
        .out2_wstrb (out2_wstrb),
        .out2_wlast (out2_wlast),
        .out2_wvalid (out2_wvalid),
        .out2_wready (out2_wready),
        .out2_bid (out2_bid),
        .out2_bresp (out2_bresp),
        .out2_bvalid (out2_bvalid),
        .out2_bready (out2_bready),
        .out2_arid (out2_arid),
        .out2_araddr (out2_araddr),
        .out2_arlen (out2_arlen),
        .out2_arsize (out2_arsize),
        .out2_arburst (out2_arburst),
        .out2_aruser (out2_aruser),
        .out2_arvalid (out2_arvalid),
        .out2_arready (out2_arready),
        .out2_rid (out2_rid),
        .out2_rdata (out2_rdata),
        .out2_rresp (out2_rresp),
        .out2_rlast (out2_rlast),
        .out2_rvalid (out2_rvalid),
        .out2_rready (out2_rready),

    `endif

    `ifdef INC_M3

        .in3_awid (in3_awid),
        .in3_awaddr (in3_awaddr),
        .in3_awlen (in3_awlen),
        .in3_awsize (in3_awsize),
        .in3_awburst (in3_awburst),
        .in3_awuser (in3_awuser),
        .in3_awvalid (in3_awvalid),
        .in3_awready (in3_awready),
        .in3_wdata (in3_wdata),
        .in3_wstrb (in3_wstrb),
        .in3_wlast (in3_wlast),
        .in3_wvalid (in3_wvalid),
        .in3_wready (in3_wready),
        .in3_bid (in3_bid),
        .in3_bresp (in3_bresp),
        .in3_bvalid (in3_bvalid),
        .in3_bready (in3_bready),
        .in3_arid (in3_arid),
        .in3_araddr (in3_araddr),
        .in3_arlen (in3_arlen),
        .in3_arsize (in3_arsize),
        .in3_arburst (in3_arburst),
        .in3_aruser (in3_aruser),
        .in3_arvalid (in3_arvalid),
        .in3_arready (in3_arready),
        .in3_rid (in3_rid),
        .in3_rdata (in3_rdata),
        .in3_rresp (in3_rresp),
        .in3_rlast (in3_rlast),
        .in3_rvalid (in3_rvalid),
        .in3_rready (in3_rready),

        .out3_awid (out3_awid),
        .out3_awaddr (out3_awaddr),
        .out3_awlen (out3_awlen),
        .out3_awsize (out3_awsize),
        .out3_awburst (out3_awburst),
        .out3_awuser (out3_awuser),
        .out3_awvalid (out3_awvalid),
        .out3_awready (out3_awready),
        .out3_wdata (out3_wdata),
        .out3_wstrb (out3_wstrb),
        .out3_wlast (out3_wlast),
        .out3_wvalid (out3_wvalid),
        .out3_wready (out3_wready),
        .out3_bid (out3_bid),
        .out3_bresp (out3_bresp),
        .out3_bvalid (out3_bvalid),
        .out3_bready (out3_bready),
        .out3_arid (out3_arid),
        .out3_araddr (out3_araddr),
        .out3_arlen (out3_arlen),
        .out3_arsize (out3_arsize),
        .out3_arburst (out3_arburst),
        .out3_aruser (out3_aruser),
        .out3_arvalid (out3_arvalid),
        .out3_arready (out3_arready),
        .out3_rid (out3_rid),
        .out3_rdata (out3_rdata),
        .out3_rresp (out3_rresp),
        .out3_rlast (out3_rlast),
        .out3_rvalid (out3_rvalid),
        .out3_rready (out3_rready),

    `endif

    `ifdef INC_M4
        .in4_awid (in4_awid),
        .in4_awaddr (in4_awaddr),
        .in4_awlen (in4_awlen),
        .in4_awsize (in4_awsize),
        .in4_awburst (in4_awburst),
        .in4_awuser (in4_awuser),
        .in4_awvalid (in4_awvalid),
        .in4_awready (in4_awready),
        .in4_wdata (in4_wdata),
        .in4_wstrb (in4_wstrb),
        .in4_wlast (in4_wlast),
        .in4_wvalid (in4_wvalid),
        .in4_wready (in4_wready),
        .in4_bid (in4_bid),
        .in4_bresp (in4_bresp),
        .in4_bvalid (in4_bvalid),
        .in4_bready (in4_bready),
        .in4_arid (in4_arid),
        .in4_araddr (in4_araddr),
        .in4_arlen (in4_arlen),
        .in4_arsize (in4_arsize),
        .in4_arburst (in4_arburst),
        .in4_aruser (in4_aruser),
        .in4_arvalid (in4_arvalid),
        .in4_arready (in4_arready),
        .in4_rid (in4_rid),
        .in4_rdata (in4_rdata),
        .in4_rresp (in4_rresp),
        .in4_rlast (in4_rlast),
        .in4_rvalid (in4_rvalid),
        .in4_rready (in4_rready),

        .out4_awid (out4_awid),
        .out4_awaddr (out4_awaddr),
        .out4_awlen (out4_awlen),
        .out4_awsize (out4_awsize),
        .out4_awburst (out4_awburst),
        .out4_awuser (out4_awuser),
        .out4_awvalid (out4_awvalid),
        .out4_awready (out4_awready),
        .out4_wdata (out4_wdata),
        .out4_wstrb (out4_wstrb),
        .out4_wlast (out4_wlast),
        .out4_wvalid (out4_wvalid),
        .out4_wready (out4_wready),
        .out4_bid (out4_bid),
        .out4_bresp (out4_bresp),
        .out4_bvalid (out4_bvalid),
        .out4_bready (out4_bready),
        .out4_arid (out4_arid),
        .out4_araddr (out4_araddr),
        .out4_arlen (out4_arlen),
        .out4_arsize (out4_arsize),
        .out4_arburst (out4_arburst),
        .out4_aruser (out4_aruser),
        .out4_arvalid (out4_arvalid),
        .out4_arready (out4_arready),
        .out4_rid (out4_rid),
        .out4_rdata (out4_rdata),
        .out4_rresp (out4_rresp),
        .out4_rlast (out4_rlast),
        .out4_rvalid (out4_rvalid),
        .out4_rready (out4_rready),

    `endif

    `ifdef INC_M5

        .in5_awid (in5_awid),
        .in5_awaddr (in5_awaddr),
        .in5_awlen (in5_awlen),
        .in5_awsize (in5_awsize),
        .in5_awburst (in5_awburst),
        .in5_awuser (in5_awuser),
        .in5_awvalid (in5_awvalid),
        .in5_awready (in5_awready),
        .in5_wdata (in5_wdata),
        .in5_wstrb (in5_wstrb),
        .in5_wlast (in5_wlast),
        .in5_wvalid (in5_wvalid),
        .in5_wready (in5_wready),
        .in5_bid (in5_bid),
        .in5_bresp (in5_bresp),
        .in5_bvalid (in5_bvalid),
        .in5_bready (in5_bready),
        .in5_arid (in5_arid),
        .in5_araddr (in5_araddr),
        .in5_arlen (in5_arlen),
        .in5_arsize (in5_arsize),
        .in5_arburst (in5_arburst),
        .in5_aruser (in5_aruser),
        .in5_arvalid (in5_arvalid),
        .in5_arready (in5_arready),
        .in5_rid (in5_rid),
        .in5_rdata (in5_rdata),
        .in5_rresp (in5_rresp),
        .in5_rlast (in5_rlast),
        .in5_rvalid (in5_rvalid),
        .in5_rready (in5_rready),

        .out5_awid (out5_awid),
        .out5_awaddr (out5_awaddr),
        .out5_awlen (out5_awlen),
        .out5_awsize (out5_awsize),
        .out5_awburst (out5_awburst),
        .out5_awuser (out5_awuser),
        .out5_awvalid (out5_awvalid),
        .out5_awready (out5_awready),
        .out5_wdata (out5_wdata),
        .out5_wstrb (out5_wstrb),
        .out5_wlast (out5_wlast),
        .out5_wvalid (out5_wvalid),
        .out5_wready (out5_wready),
        .out5_bid (out5_bid),
        .out5_bresp (out5_bresp),
        .out5_bvalid (out5_bvalid),
        .out5_bready (out5_bready),
        .out5_arid (out5_arid),
        .out5_araddr (out5_araddr),
        .out5_arlen (out5_arlen),
        .out5_arsize (out5_arsize),
        .out5_arburst (out5_arburst),
        .out5_aruser (out5_aruser),
        .out5_arvalid (out5_arvalid),
        .out5_arready (out5_arready),
        .out5_rid (out5_rid),
        .out5_rdata (out5_rdata),
        .out5_rresp (out5_rresp),
        .out5_rlast (out5_rlast),
        .out5_rvalid (out5_rvalid),
        .out5_rready (out5_rready),

    `endif

    `ifdef INC_M6

        .in6_awid (in6_awid),
        .in6_awaddr (in6_awaddr),
        .in6_awlen (in6_awlen),
        .in6_awsize (in6_awsize),
        .in6_awburst (in6_awburst),
        .in6_awuser (in6_awuser),
        .in6_awvalid (in6_awvalid),
        .in6_awready (in6_awready),
        .in6_wdata (in6_wdata),
        .in6_wstrb (in6_wstrb),
        .in6_wlast (in6_wlast),
        .in6_wvalid (in6_wvalid),
        .in6_wready (in6_wready),
        .in6_bid (in6_bid),
        .in6_bresp (in6_bresp),
        .in6_bvalid (in6_bvalid),
        .in6_bready (in6_bready),
        .in6_arid (in6_arid),
        .in6_araddr (in6_araddr),
        .in6_arlen (in6_arlen),
        .in6_arsize (in6_arsize),
        .in6_arburst (in6_arburst),
        .in6_aruser (in6_aruser),
        .in6_arvalid (in6_arvalid),
        .in6_arready (in6_arready),
        .in6_rid (in6_rid),
        .in6_rdata (in6_rdata),
        .in6_rresp (in6_rresp),
        .in6_rlast (in6_rlast),
        .in6_rvalid (in6_rvalid),
        .in6_rready (in6_rready),

        .out6_awid (out6_awid),
        .out6_awaddr (out6_awaddr),
        .out6_awlen (out6_awlen),
        .out6_awsize (out6_awsize),
        .out6_awburst (out6_awburst),
        .out6_awuser (out6_awuser),
        .out6_awvalid (out6_awvalid),
        .out6_awready (out6_awready),
        .out6_wdata (out6_wdata),
        .out6_wstrb (out6_wstrb),
        .out6_wlast (out6_wlast),
        .out6_wvalid (out6_wvalid),
        .out6_wready (out6_wready),
        .out6_bid (out6_bid),
        .out6_bresp (out6_bresp),
        .out6_bvalid (out6_bvalid),
        .out6_bready (out6_bready),
        .out6_arid (out6_arid),
        .out6_araddr (out6_araddr),
        .out6_arlen (out6_arlen),
        .out6_arsize (out6_arsize),
        .out6_arburst (out6_arburst),
        .out6_aruser (out6_aruser),
        .out6_arvalid (out6_arvalid),
        .out6_arready (out6_arready),
        .out6_rid (out6_rid),
        .out6_rdata (out6_rdata),
        .out6_rresp (out6_rresp),
        .out6_rlast (out6_rlast),
        .out6_rvalid (out6_rvalid),
        .out6_rready (out6_rready),

    `endif

    `ifdef INC_M7

        .in7_awid (in7_awid),
        .in7_awaddr (in7_awaddr),
        .in7_awlen (in7_awlen),
        .in7_awsize (in7_awsize),
        .in7_awburst (in7_awburst),
        .in7_awuser (in7_awuser),
        .in7_awvalid (in7_awvalid),
        .in7_awready (in7_awready),
        .in7_wdata (in7_wdata),
        .in7_wstrb (in7_wstrb),
        .in7_wlast (in7_wlast),
        .in7_wvalid (in7_wvalid),
        .in7_wready (in7_wready),
        .in7_bid (in7_bid),
        .in7_bresp (in7_bresp),
        .in7_bvalid (in7_bvalid),
        .in7_bready (in7_bready),
        .in7_arid (in7_arid),
        .in7_araddr (in7_araddr),
        .in7_arlen (in7_arlen),
        .in7_arsize (in7_arsize),
        .in7_arburst (in7_arburst),
        .in7_aruser (in7_aruser),
        .in7_arvalid (in7_arvalid),
        .in7_arready (in7_arready),
        .in7_rid (in7_rid),
        .in7_rdata (in7_rdata),
        .in7_rresp (in7_rresp),
        .in7_rlast (in7_rlast),
        .in7_rvalid (in7_rvalid),
        .in7_rready (in7_rready),

        .out7_awid (out7_awid),
        .out7_awaddr (out7_awaddr),
        .out7_awlen (out7_awlen),
        .out7_awsize (out7_awsize),
        .out7_awburst (out7_awburst),
        .out7_awuser (out7_awuser),
        .out7_awvalid (out7_awvalid),
        .out7_awready (out7_awready),
        .out7_wdata (out7_wdata),
        .out7_wstrb (out7_wstrb),
        .out7_wlast (out7_wlast),
        .out7_wvalid (out7_wvalid),
        .out7_wready (out7_wready),
        .out7_bid (out7_bid),
        .out7_bresp (out7_bresp),
        .out7_bvalid (out7_bvalid),
        .out7_bready (out7_bready),
        .out7_arid (out7_arid),
        .out7_araddr (out7_araddr),
        .out7_arlen (out7_arlen),
        .out7_arsize (out7_arsize),
        .out7_arburst (out7_arburst),
        .out7_aruser (out7_aruser),
        .out7_arvalid (out7_arvalid),
        .out7_arready (out7_arready),
        .out7_rid (out7_rid),
        .out7_rdata (out7_rdata),
        .out7_rresp (out7_rresp),
        .out7_rlast (out7_rlast),
        .out7_rvalid (out7_rvalid),
        .out7_rready (out7_rready),

    `endif

    `ifdef INC_M8

        .in8_awid (in8_awid),
        .in8_awaddr (in8_awaddr),
        .in8_awlen (in8_awlen),
        .in8_awsize (in8_awsize),
        .in8_awburst (in8_awburst),
        .in8_awuser (in8_awuser),
        .in8_awvalid (in8_awvalid),
        .in8_awready (in8_awready),
        .in8_wdata (in8_wdata),
        .in8_wstrb (in8_wstrb),
        .in8_wlast (in8_wlast),
        .in8_wvalid (in8_wvalid),
        .in8_wready (in8_wready),
        .in8_bid (in8_bid),
        .in8_bresp (in8_bresp),
        .in8_bvalid (in8_bvalid),
        .in8_bready (in8_bready),
        .in8_arid (in8_arid),
        .in8_araddr (in8_araddr),
        .in8_arlen (in8_arlen),
        .in8_arsize (in8_arsize),
        .in8_arburst (in8_arburst),
        .in8_aruser (in8_aruser),
        .in8_arvalid (in8_arvalid),
        .in8_arready (in8_arready),
        .in8_rid (in8_rid),
        .in8_rdata (in8_rdata),
        .in8_rresp (in8_rresp),
        .in8_rlast (in8_rlast),
        .in8_rvalid (in8_rvalid),
        .in8_rready (in8_rready),

        .out8_awid (out8_awid),
        .out8_awaddr (out8_awaddr),
        .out8_awlen (out8_awlen),
        .out8_awsize (out8_awsize),
        .out8_awburst (out8_awburst),
        .out8_awuser (out8_awuser),
        .out8_awvalid (out8_awvalid),
        .out8_awready (out8_awready),
        .out8_wdata (out8_wdata),
        .out8_wstrb (out8_wstrb),
        .out8_wlast (out8_wlast),
        .out8_wvalid (out8_wvalid),
        .out8_wready (out8_wready),
        .out8_bid (out8_bid),
        .out8_bresp (out8_bresp),
        .out8_bvalid (out8_bvalid),
        .out8_bready (out8_bready),
        .out8_arid (out8_arid),
        .out8_araddr (out8_araddr),
        .out8_arlen (out8_arlen),
        .out8_arsize (out8_arsize),
        .out8_arburst (out8_arburst),
        .out8_aruser (out8_aruser),
        .out8_arvalid (out8_arvalid),
        .out8_arready (out8_arready),
        .out8_rid (out8_rid),
        .out8_rdata (out8_rdata),
        .out8_rresp (out8_rresp),
        .out8_rlast (out8_rlast),
        .out8_rvalid (out8_rvalid),
        .out8_rready (out8_rready),

    `endif

        .bw_throt_regs (bw_throt_regs),

        .aclk (aclk),
        .aresetn (aresetn)
    );



endmodule

`default_nettype wire